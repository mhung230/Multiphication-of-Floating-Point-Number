module sum_3bits(
  